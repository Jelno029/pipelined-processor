LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

entity MEM_STAGE is
port(
		i_ctl_mem	: in std_logic_vector(2 downto 0);
		i_aluZero	: in std_logic;
		i_data		: in std_logic_vector(7 downto 0);
		i_writeData	: in std_logic_vector(7 downto 0);
		i_clk			: in std_logic;
		
		o_branchMux	: out std_logic;
		o_memData	: out std_logic_vector(7 downto 0);
		o_dataBypass: out std_logic_vector(7 downto 0));
end MEM_STAGE;


architecture mem_rtl of Mem_STAGE is

component datamem is
PORT(
		address	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		clock		: IN STD_LOGIC  := '1';
		data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		rden		: IN STD_LOGIC  := '1';
		wren		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));
end component;


begin

dmem:datamem port map(i_data, i_clk, i_writeData, i_ctl_mem(1), i_ctl_mem(0), o_memData);

o_branchMux <= i_ctl_mem(2) and i_aluZero;

end mem_rtl;